module DataPath ();
  
endmodule
