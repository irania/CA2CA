module ALUController ();
endmodule
