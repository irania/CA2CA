module ARMMicroController();
endmodule