module Controller ();
endmodule
